module vec_buffer(
    
);

endmodule